library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Filters is
	port (
		clk_i: in std_logic;
		signal_i: in integer;
		signa_o: out integer
	);
end entity;

architecture rtl of Filters is

begin

end architecture;
